`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.03.2023 20:50:35
// Design Name: 
// Module Name: mod33
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

/*
Nombre modulo: 3.3
Fecha de creaci�n: 29-03-2023
Fecha de modificaci�n: 
Funci�n: cable
*/


module cable(
    input logic A,
    output logic B
    );
    
    assign B = A;
endmodule
